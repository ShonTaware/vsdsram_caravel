VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_32_256_sky130A
   CLASS BLOCK ;
   SIZE 578.38 BY 355.34 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  131.24 0.0 131.62 1.06 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  143.48 0.0 143.86 1.06 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  157.76 0.0 158.14 1.06 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  170.0 0.0 170.38 1.06 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  182.92 0.0 183.3 1.06 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  196.52 0.0 196.9 1.06 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  209.44 0.0 209.82 1.06 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  222.36 0.0 222.74 1.06 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  235.96 0.0 236.34 1.06 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  249.56 0.0 249.94 1.06 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  262.48 0.0 262.86 1.06 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  275.4 0.0 275.78 1.06 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  288.32 0.0 288.7 1.06 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  301.24 0.0 301.62 1.06 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  314.84 0.0 315.22 1.06 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  328.44 0.0 328.82 1.06 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  340.68 0.0 341.06 1.06 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  354.28 0.0 354.66 1.06 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  367.2 0.0 367.58 1.06 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  380.8 0.0 381.18 1.06 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  393.04 0.0 393.42 1.06 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  406.64 0.0 407.02 1.06 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  420.24 0.0 420.62 1.06 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  433.16 0.0 433.54 1.06 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  445.4 0.0 445.78 1.06 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  459.0 0.0 459.38 1.06 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  471.92 0.0 472.3 1.06 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  484.84 0.0 485.22 1.06 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  499.12 0.0 499.5 1.06 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  512.04 0.0 512.42 1.06 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  524.28 0.0 524.66 1.06 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  537.88 0.0 538.26 1.06 ;
      END
   END din0[31]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  104.72 0.0 105.1 1.06 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  117.64 0.0 118.02 1.06 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 132.6 1.06 132.98 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 135.32 1.06 135.7 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 141.44 1.06 141.82 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 143.48 1.06 143.86 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 150.28 1.06 150.66 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 151.64 1.06 152.02 ;
      END
   END addr0[7]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 20.4 1.06 20.78 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 22.44 1.06 22.82 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  38.08 0.0 38.46 1.06 ;
      END
   END clk0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  140.76 0.0 141.14 1.06 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  153.68 0.0 154.06 1.06 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  166.6 0.0 166.98 1.06 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  179.52 0.0 179.9 1.06 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  193.12 0.0 193.5 1.06 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  206.04 0.0 206.42 1.06 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  218.96 0.0 219.34 1.06 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  232.56 0.0 232.94 1.06 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  245.48 0.0 245.86 1.06 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  258.4 0.0 258.78 1.06 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  272.0 0.0 272.38 1.06 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  284.92 0.0 285.3 1.06 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  297.84 0.0 298.22 1.06 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  311.44 0.0 311.82 1.06 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  324.36 0.0 324.74 1.06 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  337.28 0.0 337.66 1.06 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  350.88 0.0 351.26 1.06 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  363.8 0.0 364.18 1.06 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  377.4 0.0 377.78 1.06 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  391.0 0.0 391.38 1.06 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  403.24 0.0 403.62 1.06 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  417.52 0.0 417.9 1.06 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  430.44 0.0 430.82 1.06 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  443.36 0.0 443.74 1.06 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  456.28 0.0 456.66 1.06 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  469.2 0.0 469.58 1.06 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  482.8 0.0 483.18 1.06 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  495.72 0.0 496.1 1.06 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  509.32 0.0 509.7 1.06 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  522.24 0.0 522.62 1.06 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  535.16 0.0 535.54 1.06 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  577.32 33.32 578.38 33.7 ;
      END
   END dout0[31]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  4.76 4.76 6.5 351.94 ;
         LAYER met3 ;
         RECT  4.76 4.76 573.62 6.5 ;
         LAYER met3 ;
         RECT  4.76 350.2 573.62 351.94 ;
         LAYER met4 ;
         RECT  571.88 4.76 573.62 351.94 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  575.28 1.36 577.02 355.34 ;
         LAYER met3 ;
         RECT  1.36 353.6 577.02 355.34 ;
         LAYER met3 ;
         RECT  1.36 1.36 577.02 3.1 ;
         LAYER met4 ;
         RECT  1.36 1.36 3.1 355.34 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 577.76 354.72 ;
   LAYER  met2 ;
      RECT  0.62 0.62 577.76 354.72 ;
   LAYER  met3 ;
      RECT  1.66 132.0 577.76 133.58 ;
      RECT  0.62 133.58 1.66 134.72 ;
      RECT  0.62 136.3 1.66 140.84 ;
      RECT  0.62 142.42 1.66 142.88 ;
      RECT  0.62 144.46 1.66 149.68 ;
      RECT  0.62 21.38 1.66 21.84 ;
      RECT  0.62 23.42 1.66 132.0 ;
      RECT  1.66 32.72 576.72 34.3 ;
      RECT  1.66 34.3 576.72 132.0 ;
      RECT  576.72 34.3 577.76 132.0 ;
      RECT  1.66 4.16 4.16 7.1 ;
      RECT  1.66 7.1 4.16 32.72 ;
      RECT  4.16 7.1 574.22 32.72 ;
      RECT  574.22 4.16 576.72 7.1 ;
      RECT  574.22 7.1 576.72 32.72 ;
      RECT  1.66 133.58 4.16 349.6 ;
      RECT  1.66 349.6 4.16 352.54 ;
      RECT  4.16 133.58 574.22 349.6 ;
      RECT  574.22 133.58 577.76 349.6 ;
      RECT  574.22 349.6 577.76 352.54 ;
      RECT  0.62 152.62 0.76 353.0 ;
      RECT  0.62 353.0 0.76 354.72 ;
      RECT  0.76 152.62 1.66 353.0 ;
      RECT  1.66 352.54 4.16 353.0 ;
      RECT  4.16 352.54 574.22 353.0 ;
      RECT  574.22 352.54 577.62 353.0 ;
      RECT  577.62 352.54 577.76 353.0 ;
      RECT  577.62 353.0 577.76 354.72 ;
      RECT  0.62 0.62 0.76 0.76 ;
      RECT  0.62 0.76 0.76 3.7 ;
      RECT  0.62 3.7 0.76 19.8 ;
      RECT  0.76 0.62 1.66 0.76 ;
      RECT  0.76 3.7 1.66 19.8 ;
      RECT  576.72 0.62 577.62 0.76 ;
      RECT  576.72 3.7 577.62 32.72 ;
      RECT  577.62 0.62 577.76 0.76 ;
      RECT  577.62 0.76 577.76 3.7 ;
      RECT  577.62 3.7 577.76 32.72 ;
      RECT  1.66 0.62 4.16 0.76 ;
      RECT  1.66 3.7 4.16 4.16 ;
      RECT  4.16 0.62 574.22 0.76 ;
      RECT  4.16 3.7 574.22 4.16 ;
      RECT  574.22 0.62 576.72 0.76 ;
      RECT  574.22 3.7 576.72 4.16 ;
   LAYER  met4 ;
      RECT  130.64 1.66 132.22 354.72 ;
      RECT  105.7 0.62 117.04 1.66 ;
      RECT  118.62 0.62 130.64 1.66 ;
      RECT  39.06 0.62 104.12 1.66 ;
      RECT  132.22 0.62 140.16 1.66 ;
      RECT  141.74 0.62 142.88 1.66 ;
      RECT  144.46 0.62 153.08 1.66 ;
      RECT  154.66 0.62 157.16 1.66 ;
      RECT  158.74 0.62 166.0 1.66 ;
      RECT  167.58 0.62 169.4 1.66 ;
      RECT  170.98 0.62 178.92 1.66 ;
      RECT  180.5 0.62 182.32 1.66 ;
      RECT  183.9 0.62 192.52 1.66 ;
      RECT  194.1 0.62 195.92 1.66 ;
      RECT  197.5 0.62 205.44 1.66 ;
      RECT  207.02 0.62 208.84 1.66 ;
      RECT  210.42 0.62 218.36 1.66 ;
      RECT  219.94 0.62 221.76 1.66 ;
      RECT  223.34 0.62 231.96 1.66 ;
      RECT  233.54 0.62 235.36 1.66 ;
      RECT  236.94 0.62 244.88 1.66 ;
      RECT  246.46 0.62 248.96 1.66 ;
      RECT  250.54 0.62 257.8 1.66 ;
      RECT  259.38 0.62 261.88 1.66 ;
      RECT  263.46 0.62 271.4 1.66 ;
      RECT  272.98 0.62 274.8 1.66 ;
      RECT  276.38 0.62 284.32 1.66 ;
      RECT  285.9 0.62 287.72 1.66 ;
      RECT  289.3 0.62 297.24 1.66 ;
      RECT  298.82 0.62 300.64 1.66 ;
      RECT  302.22 0.62 310.84 1.66 ;
      RECT  312.42 0.62 314.24 1.66 ;
      RECT  315.82 0.62 323.76 1.66 ;
      RECT  325.34 0.62 327.84 1.66 ;
      RECT  329.42 0.62 336.68 1.66 ;
      RECT  338.26 0.62 340.08 1.66 ;
      RECT  341.66 0.62 350.28 1.66 ;
      RECT  351.86 0.62 353.68 1.66 ;
      RECT  355.26 0.62 363.2 1.66 ;
      RECT  364.78 0.62 366.6 1.66 ;
      RECT  368.18 0.62 376.8 1.66 ;
      RECT  378.38 0.62 380.2 1.66 ;
      RECT  381.78 0.62 390.4 1.66 ;
      RECT  391.98 0.62 392.44 1.66 ;
      RECT  394.02 0.62 402.64 1.66 ;
      RECT  404.22 0.62 406.04 1.66 ;
      RECT  407.62 0.62 416.92 1.66 ;
      RECT  418.5 0.62 419.64 1.66 ;
      RECT  421.22 0.62 429.84 1.66 ;
      RECT  431.42 0.62 432.56 1.66 ;
      RECT  434.14 0.62 442.76 1.66 ;
      RECT  444.34 0.62 444.8 1.66 ;
      RECT  446.38 0.62 455.68 1.66 ;
      RECT  457.26 0.62 458.4 1.66 ;
      RECT  459.98 0.62 468.6 1.66 ;
      RECT  470.18 0.62 471.32 1.66 ;
      RECT  472.9 0.62 482.2 1.66 ;
      RECT  483.78 0.62 484.24 1.66 ;
      RECT  485.82 0.62 495.12 1.66 ;
      RECT  496.7 0.62 498.52 1.66 ;
      RECT  500.1 0.62 508.72 1.66 ;
      RECT  510.3 0.62 511.44 1.66 ;
      RECT  513.02 0.62 521.64 1.66 ;
      RECT  523.22 0.62 523.68 1.66 ;
      RECT  525.26 0.62 534.56 1.66 ;
      RECT  536.14 0.62 537.28 1.66 ;
      RECT  4.16 1.66 7.1 4.16 ;
      RECT  4.16 352.54 7.1 354.72 ;
      RECT  7.1 1.66 130.64 4.16 ;
      RECT  7.1 4.16 130.64 352.54 ;
      RECT  7.1 352.54 130.64 354.72 ;
      RECT  132.22 1.66 571.28 4.16 ;
      RECT  132.22 4.16 571.28 352.54 ;
      RECT  132.22 352.54 571.28 354.72 ;
      RECT  571.28 1.66 574.22 4.16 ;
      RECT  571.28 352.54 574.22 354.72 ;
      RECT  538.86 0.62 574.68 0.76 ;
      RECT  538.86 0.76 574.68 1.66 ;
      RECT  574.68 0.62 577.62 0.76 ;
      RECT  577.62 0.62 577.76 0.76 ;
      RECT  577.62 0.76 577.76 1.66 ;
      RECT  574.22 1.66 574.68 4.16 ;
      RECT  577.62 1.66 577.76 4.16 ;
      RECT  574.22 4.16 574.68 352.54 ;
      RECT  577.62 4.16 577.76 352.54 ;
      RECT  574.22 352.54 574.68 354.72 ;
      RECT  577.62 352.54 577.76 354.72 ;
      RECT  0.62 0.62 0.76 0.76 ;
      RECT  0.62 0.76 0.76 1.66 ;
      RECT  0.76 0.62 3.7 0.76 ;
      RECT  3.7 0.62 37.48 0.76 ;
      RECT  3.7 0.76 37.48 1.66 ;
      RECT  0.62 1.66 0.76 4.16 ;
      RECT  3.7 1.66 4.16 4.16 ;
      RECT  0.62 4.16 0.76 352.54 ;
      RECT  3.7 4.16 4.16 352.54 ;
      RECT  0.62 352.54 0.76 354.72 ;
      RECT  3.7 352.54 4.16 354.72 ;
   END
END    sram_32_256_sky130A
END    LIBRARY
