* SPICE3 file created from sky130_vsdinv_1x.ext - technology: sky130A

.subckt pinv
X0 Z A gnd gnd sky130_fd_pr__nfet_01v8 w=43 l=15
X1 Z A vdd vdd sky130_fd_pr__pfet_01v8 w=70 l=15


.ends
