.subckt pnand2
X0 NET1 A Z gnd sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u
X1 NET1 B gnd gnd sky130_fd_pr__nfet_01v8 w=0.42u l=0.15u

X2 Z A vdd vdd sky130_fd_pr__pfet_01v8 w=0.97u l=0.15u
X3 Z B vdd vdd sky130_fd_pr__pfet_01v8 w=0.97u l=0.15u
.ends
